module pps (clk1,clk2);
input   clk1;
output  wire clk2;

assign clk2=clk1;


endmodule