module ten (ten1,ten2);
input   ten1;
output  wire ten2;

assign ten2=ten1;


endmodule