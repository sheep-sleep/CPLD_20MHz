module transmit_en(transmit_en1,transmit_en2);
input   transmit_en1;
output  wire transmit_en2;

assign transmit_en2=transmit_en1;

endmodule